
//=======================================================
//  MODULE Definition
//=======================================================

module SC_STATEMACHINE_ENVIRONMENT 
(
	//////////// INPUTS //////////
	SC_STATEMACHINE_ENVIRONMENT_CLOCK_50,
	SC_STATEMACHINE_ENVIRONMENT_RESET_InLow,
	SC_STATEMACHINE_ENVIRONMENT_START_InLow,
	SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow,	
	SC_STATEMACHINE_ENVIRONMENT_LOSE_InLow,
	SC_STATEMACHINE_ENVIRONMENT_WIN_InLow,
	SC_STATEMACHINE_ENVIRONMENT_DOWN_InLow,
	SC_STATEMACHINE_ENVIRONMENT_LEVEL_InBus,
	
	//////////// OUTPUTS //////////
	SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out,
	SC_STATEMACHINE_ENVIRONMENT_LOAD_Out,
	SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out,
	SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out,
	SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus
);	

//=======================================================
//  PARAMETER declarations
//=======================================================

localparam STATE_RESET									= 0;
localparam STATE_START									= 1;
localparam STATE_TRANSITION							= 2;
localparam STATE_READY1									= 4;
localparam STATE_READY2									= 12;
localparam STATE_READY3									= 13;
localparam STATE_SHIFTDOWN_0							= 5; 
localparam STATE_SHIFTDOWN_1							= 6;
localparam STATE_SHIFTDOWN_02							= 14; 
localparam STATE_SHIFTDOWN_12							= 15;
localparam STATE_SHIFTDOWN_03							= 16; 
localparam STATE_SHIFTDOWN_13							= 17;
localparam STATE_LOSE									= 7;	
localparam STATE_WIN										= 8;
localparam STATE_TRANSITION1							= 9;
localparam STATE_TRANSITION2							= 10;
localparam STATE_TRANSITION3							= 11;

//=======================================================
//  PORT declarations
//=======================================================

input	SC_STATEMACHINE_ENVIRONMENT_CLOCK_50;
input	SC_STATEMACHINE_ENVIRONMENT_RESET_InLow;
input	SC_STATEMACHINE_ENVIRONMENT_START_InLow;
input	SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow;	
input	SC_STATEMACHINE_ENVIRONMENT_LOSE_InLow;
input	SC_STATEMACHINE_ENVIRONMENT_WIN_InLow;
input SC_STATEMACHINE_ENVIRONMENT_DOWN_InLow;
input[2:0] SC_STATEMACHINE_ENVIRONMENT_LEVEL_InBus;
	
output reg	SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out;
output reg	SC_STATEMACHINE_ENVIRONMENT_LOAD_Out;
output reg  SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out;
output reg	SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out;
output reg[2:0]	SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus;

//=======================================================
//  REG/WIRE declarations
//=======================================================
reg [7:0] STATE_Register;
reg [7:0] STATE_Signal;
//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
// NEXT STATE LOGIC : COMBINATIONAL
always @(*)
begin
	case (STATE_Register)
		
		STATE_RESET: 	STATE_Signal = STATE_START;
		
		STATE_START: 	if (SC_STATEMACHINE_ENVIRONMENT_START_InLow == 1'b0) 
								STATE_Signal = STATE_TRANSITION;
							else 
								STATE_Signal = STATE_START;
								
		STATE_TRANSITION: if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
									STATE_Signal = STATE_TRANSITION1;
								else 
									STATE_Signal = STATE_TRANSITION;
									
		STATE_TRANSITION1: if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
									STATE_Signal = STATE_READY1;
								else 
									STATE_Signal = STATE_TRANSITION1;
								
		STATE_READY1: if (SC_STATEMACHINE_ENVIRONMENT_LEVEL_InBus == 2'b10)
							 STATE_Signal = STATE_TRANSITION2; 
						 else if (SC_STATEMACHINE_ENVIRONMENT_LOSE_InLow == 1'b0)
							 STATE_Signal = STATE_LOSE;
						 else if (SC_STATEMACHINE_ENVIRONMENT_WIN_InLow == 1'b0)
						    STATE_Signal = STATE_WIN;
						 else if (SC_STATEMACHINE_ENVIRONMENT_DOWN_InLow == 1'b0)
							 STATE_Signal = STATE_SHIFTDOWN_0;
						 else
							 STATE_Signal = STATE_READY1;
							 
		STATE_TRANSITION2: if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
									STATE_Signal = STATE_READY2;
								 else 
									STATE_Signal = STATE_TRANSITION2;
									
		STATE_READY2: if (SC_STATEMACHINE_ENVIRONMENT_LEVEL_InBus == 2'b11)
							 STATE_Signal = STATE_TRANSITION3;
						 else if (SC_STATEMACHINE_ENVIRONMENT_LOSE_InLow == 1'b0)
							 STATE_Signal = STATE_LOSE;
						 else if (SC_STATEMACHINE_ENVIRONMENT_WIN_InLow == 1'b0)
						    STATE_Signal = STATE_WIN;
						 else if (SC_STATEMACHINE_ENVIRONMENT_DOWN_InLow == 1'b0)
							 STATE_Signal = STATE_SHIFTDOWN_02;
						 else
							 STATE_Signal = STATE_READY2;
								
		STATE_TRANSITION3: if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
									STATE_Signal = STATE_READY3;
								else 
									STATE_Signal = STATE_TRANSITION3;
									
		STATE_READY3: if (SC_STATEMACHINE_ENVIRONMENT_LOSE_InLow == 1'b0)
							 STATE_Signal = STATE_LOSE;
						 else if (SC_STATEMACHINE_ENVIRONMENT_WIN_InLow == 1'b0)
						    STATE_Signal = STATE_WIN;
						 else if (SC_STATEMACHINE_ENVIRONMENT_DOWN_InLow == 1'b0)
							 STATE_Signal = STATE_SHIFTDOWN_03;
						 else
							 STATE_Signal = STATE_READY3;
		
		STATE_SHIFTDOWN_0: 	STATE_Signal = STATE_SHIFTDOWN_1;
		
		STATE_SHIFTDOWN_1: 	STATE_Signal = STATE_READY1;
		
		STATE_SHIFTDOWN_02: 	STATE_Signal = STATE_SHIFTDOWN_12;
		
		STATE_SHIFTDOWN_12: 	STATE_Signal = STATE_READY2;
		
		STATE_SHIFTDOWN_03: 	STATE_Signal = STATE_SHIFTDOWN_13;
		
		STATE_SHIFTDOWN_13: 	STATE_Signal = STATE_READY3;
		
		STATE_LOSE: if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
							STATE_Signal = STATE_RESET;
						else 
							STATE_Signal = STATE_LOSE;
		
		STATE_WIN: 	if (SC_STATEMACHINE_ENVIRONMENT_TRANSITION_InLow == 1'b0) 
							STATE_Signal = STATE_RESET;
						else 
							STATE_Signal = STATE_WIN;
		
		default : STATE_Signal = STATE_RESET;
	
	endcase
end
// STATE REGISTER : SEQUENTIAL
always @ ( posedge SC_STATEMACHINE_ENVIRONMENT_CLOCK_50 , negedge SC_STATEMACHINE_ENVIRONMENT_RESET_InLow)
begin
	if (SC_STATEMACHINE_ENVIRONMENT_RESET_InLow == 1'b0)
		STATE_Register <= STATE_RESET;
	else
		STATE_Register <= STATE_Signal;
end
//=======================================================
//  Outputs
//=======================================================
// OUTPUT LOGIC : COMBINATIONAL
always @ (*)
begin
	case (STATE_Register)
		
		STATE_RESET:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_START:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end			
								
		STATE_TRANSITION: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b001;	
		end
		
		STATE_TRANSITION1: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b100;	
		end
		
		STATE_TRANSITION2: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b101;	
		end
		
		STATE_TRANSITION3: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b110;	
		end
		
		STATE_READY1:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_READY2:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_READY3:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_0: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_1: 	
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_02: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_12: 	
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_03: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_SHIFTDOWN_13: 	
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
		
		STATE_LOSE: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b010;	
		end
		
		STATE_WIN: 
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b0;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b011;	
		end
		
		default:
		begin
			SC_STATEMACHINE_ENVIRONMENT_CLEAR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_LOAD_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_ENABLECOUNT_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SCREENSELECTOR_Out = 1'b1;
			SC_STATEMACHINE_ENVIRONMENT_SELECTIONTRAN_OutBus = 3'b000;	
		end
	endcase
end
endmodule
