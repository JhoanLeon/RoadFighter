
//=======================================================
//  MODULE Definition
//=======================================================

module SC_REGISTER_ENVIRONMENT
(

//////////// INPUTS //////////
SC_REGISTER_ENVIRONMENT_CLOCK_50,
SC_REGISTER_ENVIRONMENT_RESET_InLow,
SC_REGISTER_ENVIRONMENT_clear_InLow, 
SC_REGISTER_ENVIRONMENT_load_InLow, 
SC_REGISTER_ENVIRONMENT_data_InBUS,
	
//////////// OUTPUTS //////////
SC_REGISTER_ENVIRONMENT_data7_OutBUS,
SC_REGISTER_ENVIRONMENT_data6_OutBUS,
SC_REGISTER_ENVIRONMENT_data5_OutBUS,
SC_REGISTER_ENVIRONMENT_data4_OutBUS,
SC_REGISTER_ENVIRONMENT_data3_OutBUS,
SC_REGISTER_ENVIRONMENT_data2_OutBUS,
SC_REGISTER_ENVIRONMENT_data1_OutBUS,
SC_REGISTER_ENVIRONMENT_data0_OutBUS

);

//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
input		SC_REGISTER_ENVIRONMENT_CLOCK_50;
input		SC_REGISTER_ENVIRONMENT_RESET_InLow;
input		SC_REGISTER_ENVIRONMENT_clear_InLow;
input		SC_REGISTER_ENVIRONMENT_load_InLow;	
input		[7:0]	SC_REGISTER_ENVIRONMENT_data_InBUS;

output wire[7:0]	SC_REGISTER_ENVIRONMENT_data7_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data6_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data5_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data4_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data3_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data2_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data1_OutBUS;
output wire[7:0]	SC_REGISTER_ENVIRONMENT_data0_OutBUS;

//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================

SC_REGGENERAL SC_REGGENERAL_u7 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data_InBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data7_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u6 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data7_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data6_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u5 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data6_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data5_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u4 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data5_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data4_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u3 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data4_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data3_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u2 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data3_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data2_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u1 
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data2_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data1_OutBUS)

);

SC_REGGENERAL SC_REGGENERAL_u0
(

.SC_REGGENERAL_CLOCK_50(SC_REGISTER_ENVIRONMENT_CLOCK_50),
.SC_REGGENERAL_RESET_InLow(SC_REGISTER_ENVIRONMENT_RESET_InLow),
.SC_REGGENERAL_clear_InLow(SC_REGISTER_ENVIRONMENT_clear_InLow), 
.SC_REGGENERAL_load_InLow(SC_REGISTER_ENVIRONMENT_load_InLow), 
.SC_REGGENERAL_data_InBUS(SC_REGISTER_ENVIRONMENT_data1_OutBUS),
	
.SC_REGGENERAL_data_OutBUS(SC_REGISTER_ENVIRONMENT_data0_OutBUS)

);

endmodule
